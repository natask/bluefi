//----------------------------------------------------------------------//
// The MIT License 
// 
// Copyright (c) 2007 Alfred Man Cheuk Ng, mcn02@mit.edu 
// 
// Permission is hereby granted, free of charge, to any person 
// obtaining a copy of this software and associated documentation 
// files (the "Software"), to deal in the Software without 
// restriction, including without limitation the rights to use,
// copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
// OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
// HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
// WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
// FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
// OTHER DEALINGS IN THE SOFTWARE.
//----------------------------------------------------------------------//

import BRAMFIFO::*;
import FIFO::*;

(* synthesize *)
module mkBRAMFIFOTest (Empty);
   
   // constants
   Bit#(1) lo_index = 0;
   Bit#(1) hi_index = 1;
   
   // state elements
   Reg#(Bit#(32)) cycle <- mkReg(0);
   FIFO#(Bit#(32)) fifo <- mkBRAMFIFO(lo_index,hi_index);
   
   // rules
   rule enqFIFO (True);
      fifo.enq(cycle);
      $display("Enq data: %d at cycle %d", cycle, cycle);
   endrule
   
   rule readFIFO (True);
      $display("First data: %d at cycle %d", fifo.first, cycle);
   endrule
   
   rule deqFIFO (cycle[1:0] == 0);
      fifo.deq();
      $display("Deq data: %d at cycle %d", fifo.first, cycle);
   endrule
   
   rule tick (True);
      cycle <= cycle + 1;
      if (cycle == 100000)
	 $finish;
   endrule   
endmodule