//----------------------------------------------------------------------//
// The MIT License 
// 
// Copyright (c) 2007 Alfred Man Cheuk Ng, mcn02@mit.edu 
// 
// Permission is hereby granted, free of charge, to any person 
// obtaining a copy of this software and associated documentation 
// files (the "Software"), to deal in the Software without 
// restriction, including without limitation the rights to use,
// copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
// OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
// HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
// WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
// FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
// OTHER DEALINGS IN THE SOFTWARE.
//----------------------------------------------------------------------//

import List::*;
import Vector::*;
import Complex::*;
import DataTypes::*;
import RegFile::*;
import FixedPoint::*;
import FPComplex::*;

// function to generate short training sequence
function Vector#(256, FPComplex#(2,14)) getShortPreambles();
	Vector#(256, FPComplex#(2,14)) tempV = Vector::toVector(
		List::cons(cmplx(fromRational(625000,10000000), fromRational(625000,10000000)),
		List::cons(cmplx(fromRational(353100,10000000), fromRational(-1029300,10000000)),
		List::cons(cmplx(fromRational(-757100,10000000), fromRational(194400,10000000)),
		List::cons(cmplx(fromRational(-441500,10000000), fromRational(665000,10000000)),
		List::cons(cmplx(fromRational(369300,10000000), fromRational(-62800,10000000)),
		List::cons(cmplx(fromRational(920500,10000000), fromRational(597200,10000000)),
		List::cons(cmplx(fromRational(347100,10000000), fromRational(-294900,10000000)),
		List::cons(cmplx(fromRational(206500,10000000), fromRational(-921400,10000000)),
		List::cons(cmplx(fromRational(552400,10000000), fromRational(-552400,10000000)),
		List::cons(cmplx(fromRational(-10100,10000000), fromRational(-169700,10000000)),
		List::cons(cmplx(fromRational(-34800,10000000), fromRational(558900,10000000)),
		List::cons(cmplx(fromRational(-239100,10000000), fromRational(-507500,10000000)),
		List::cons(cmplx(fromRational(-1021400,10000000), fromRational(-284700,10000000)),
		List::cons(cmplx(fromRational(-312000,10000000), fromRational(869900,10000000)),
		List::cons(cmplx(fromRational(766700,10000000), fromRational(-538200,10000000)),
		List::cons(cmplx(fromRational(-103800,10000000), fromRational(-519300,10000000)),
		List::cons(cmplx(fromRational(-1093800,10000000), fromRational(-156200,10000000)),
		List::cons(cmplx(fromRational(-160700,10000000), fromRational(-690600,10000000)),
		List::cons(cmplx(fromRational(-77700,10000000), fromRational(508300,10000000)),
		List::cons(cmplx(fromRational(-821800,10000000), fromRational(383000,10000000)),
		List::cons(cmplx(fromRational(-21700,10000000), fromRational(-623000,10000000)),
		List::cons(cmplx(fromRational(576500,10000000), fromRational(-112100,10000000)),
		List::cons(cmplx(fromRational(889200,10000000), fromRational(406700,10000000)),
		List::cons(cmplx(fromRational(400100,10000000), fromRational(645400,10000000)),
		List::cons(cmplx(fromRational(-773400,10000000), fromRational(773400,10000000)),
		List::cons(cmplx(fromRational(303000,10000000), fromRational(789100,10000000)),
		List::cons(cmplx(fromRational(471400,10000000), fromRational(-193200,10000000)),
		List::cons(cmplx(fromRational(-805300,10000000), fromRational(-747500,10000000)),
		List::cons(cmplx(fromRational(-359400,10000000), fromRational(753800,10000000)),
		List::cons(cmplx(fromRational(-303100,10000000), fromRational(727700,10000000)),
		List::cons(cmplx(fromRational(127500,10000000), fromRational(-13700,10000000)),
		List::cons(cmplx(fromRational(876900,10000000), fromRational(655200,10000000)),
		List::cons(cmplx(fromRational(0,10000000), fromRational(0,10000000)),
		List::cons(cmplx(fromRational(81500,10000000), fromRational(-850300,10000000)),
		List::cons(cmplx(fromRational(775300,10000000), fromRational(-753700,10000000)),
		List::cons(cmplx(fromRational(875700,10000000), fromRational(-480000,10000000)),
		List::cons(cmplx(fromRational(827100,10000000), fromRational(634200,10000000)),
		List::cons(cmplx(fromRational(328700,10000000), fromRational(629200,10000000)),
		List::cons(cmplx(fromRational(259700,10000000), fromRational(-300800,10000000)),
		List::cons(cmplx(fromRational(-244500,10000000), fromRational(337300,10000000)),
		List::cons(cmplx(fromRational(-552400,10000000), fromRational(552400,10000000)),
		List::cons(cmplx(fromRational(718800,10000000), fromRational(-143500,10000000)),
		List::cons(cmplx(fromRational(833200,10000000), fromRational(478600,10000000)),
		List::cons(cmplx(fromRational(-129400,10000000), fromRational(371600,10000000)),
		List::cons(cmplx(fromRational(83900,10000000), fromRational(-911700,10000000)),
		List::cons(cmplx(fromRational(598800,10000000), fromRational(-279400,10000000)),
		List::cons(cmplx(fromRational(214700,10000000), fromRational(655500,10000000)),
		List::cons(cmplx(fromRational(-439100,10000000), fromRational(678400,10000000)),
		List::cons(cmplx(fromRational(-781200,10000000), fromRational(781200,10000000)),
		List::cons(cmplx(fromRational(-1006600,10000000), fromRational(-149600,10000000)),
		List::cons(cmplx(fromRational(-382500,10000000), fromRational(-391000,10000000)),
		List::cons(cmplx(fromRational(-101900,10000000), fromRational(45900,10000000)),
		List::cons(cmplx(fromRational(-549600,10000000), fromRational(-573400,10000000)),
		List::cons(cmplx(fromRational(296900,10000000), fromRational(112400,10000000)),
		List::cons(cmplx(fromRational(195900,10000000), fromRational(630800,10000000)),
		List::cons(cmplx(fromRational(-306100,10000000), fromRational(-535100,10000000)),
		List::cons(cmplx(fromRational(773400,10000000), fromRational(-773400,10000000)),
		List::cons(cmplx(fromRational(87100,10000000), fromRational(-407700,10000000)),
		List::cons(cmplx(fromRational(-827800,10000000), fromRational(-402500,10000000)),
		List::cons(cmplx(fromRational(-470600,10000000), fromRational(-614400,10000000)),
		List::cons(cmplx(fromRational(-578100,10000000), fromRational(-182400,10000000)),
		List::cons(cmplx(fromRational(27400,10000000), fromRational(106700,10000000)),
		List::cons(cmplx(fromRational(-300900,10000000), fromRational(-545500,10000000)),
		List::cons(cmplx(fromRational(-756300,10000000), fromRational(543200,10000000)),
		List::cons(cmplx(fromRational(625000,10000000), fromRational(625000,10000000)),
		List::cons(cmplx(fromRational(353100,10000000), fromRational(-1029300,10000000)),
		List::cons(cmplx(fromRational(-757100,10000000), fromRational(194400,10000000)),
		List::cons(cmplx(fromRational(-441500,10000000), fromRational(665000,10000000)),
		List::cons(cmplx(fromRational(369300,10000000), fromRational(-62800,10000000)),
		List::cons(cmplx(fromRational(920500,10000000), fromRational(597200,10000000)),
		List::cons(cmplx(fromRational(347100,10000000), fromRational(-294900,10000000)),
		List::cons(cmplx(fromRational(206500,10000000), fromRational(-921400,10000000)),
		List::cons(cmplx(fromRational(552400,10000000), fromRational(-552400,10000000)),
		List::cons(cmplx(fromRational(-10100,10000000), fromRational(-169700,10000000)),
		List::cons(cmplx(fromRational(-34800,10000000), fromRational(558900,10000000)),
		List::cons(cmplx(fromRational(-239100,10000000), fromRational(-507500,10000000)),
		List::cons(cmplx(fromRational(-1021400,10000000), fromRational(-284700,10000000)),
		List::cons(cmplx(fromRational(-312000,10000000), fromRational(869900,10000000)),
		List::cons(cmplx(fromRational(766700,10000000), fromRational(-538200,10000000)),
		List::cons(cmplx(fromRational(-103800,10000000), fromRational(-519300,10000000)),
		List::cons(cmplx(fromRational(-1093800,10000000), fromRational(-156200,10000000)),
		List::cons(cmplx(fromRational(-160700,10000000), fromRational(-690600,10000000)),
		List::cons(cmplx(fromRational(-77700,10000000), fromRational(508300,10000000)),
		List::cons(cmplx(fromRational(-821800,10000000), fromRational(383000,10000000)),
		List::cons(cmplx(fromRational(-21700,10000000), fromRational(-623000,10000000)),
		List::cons(cmplx(fromRational(576500,10000000), fromRational(-112100,10000000)),
		List::cons(cmplx(fromRational(889200,10000000), fromRational(406700,10000000)),
		List::cons(cmplx(fromRational(400100,10000000), fromRational(645400,10000000)),
		List::cons(cmplx(fromRational(-773400,10000000), fromRational(773400,10000000)),
		List::cons(cmplx(fromRational(303000,10000000), fromRational(789100,10000000)),
		List::cons(cmplx(fromRational(471400,10000000), fromRational(-193200,10000000)),
		List::cons(cmplx(fromRational(-805300,10000000), fromRational(-747500,10000000)),
		List::cons(cmplx(fromRational(-359400,10000000), fromRational(753800,10000000)),
		List::cons(cmplx(fromRational(-303100,10000000), fromRational(727700,10000000)),
		List::cons(cmplx(fromRational(127500,10000000), fromRational(-13700,10000000)),
		List::cons(cmplx(fromRational(876900,10000000), fromRational(655200,10000000)),
		List::cons(cmplx(fromRational(0,10000000), fromRational(0,10000000)),
		List::cons(cmplx(fromRational(81500,10000000), fromRational(-850300,10000000)),
		List::cons(cmplx(fromRational(775300,10000000), fromRational(-753700,10000000)),
		List::cons(cmplx(fromRational(875700,10000000), fromRational(-480000,10000000)),
		List::cons(cmplx(fromRational(827100,10000000), fromRational(634200,10000000)),
		List::cons(cmplx(fromRational(328700,10000000), fromRational(629200,10000000)),
		List::cons(cmplx(fromRational(259700,10000000), fromRational(-300800,10000000)),
		List::cons(cmplx(fromRational(-244500,10000000), fromRational(337300,10000000)),
		List::cons(cmplx(fromRational(-552400,10000000), fromRational(552400,10000000)),
		List::cons(cmplx(fromRational(718800,10000000), fromRational(-143500,10000000)),
		List::cons(cmplx(fromRational(833200,10000000), fromRational(478600,10000000)),
		List::cons(cmplx(fromRational(-129400,10000000), fromRational(371600,10000000)),
		List::cons(cmplx(fromRational(83900,10000000), fromRational(-911700,10000000)),
		List::cons(cmplx(fromRational(598800,10000000), fromRational(-279400,10000000)),
		List::cons(cmplx(fromRational(214700,10000000), fromRational(655500,10000000)),
		List::cons(cmplx(fromRational(-439100,10000000), fromRational(678400,10000000)),
		List::cons(cmplx(fromRational(-781200,10000000), fromRational(781200,10000000)),
		List::cons(cmplx(fromRational(-1006600,10000000), fromRational(-149600,10000000)),
		List::cons(cmplx(fromRational(-382500,10000000), fromRational(-391000,10000000)),
		List::cons(cmplx(fromRational(-101900,10000000), fromRational(45900,10000000)),
		List::cons(cmplx(fromRational(-549600,10000000), fromRational(-573400,10000000)),
		List::cons(cmplx(fromRational(296900,10000000), fromRational(112400,10000000)),
		List::cons(cmplx(fromRational(195900,10000000), fromRational(630800,10000000)),
		List::cons(cmplx(fromRational(-306100,10000000), fromRational(-535100,10000000)),
		List::cons(cmplx(fromRational(773400,10000000), fromRational(-773400,10000000)),
		List::cons(cmplx(fromRational(87100,10000000), fromRational(-407700,10000000)),
		List::cons(cmplx(fromRational(-827800,10000000), fromRational(-402500,10000000)),
		List::cons(cmplx(fromRational(-470600,10000000), fromRational(-614400,10000000)),
		List::cons(cmplx(fromRational(-578100,10000000), fromRational(-182400,10000000)),
		List::cons(cmplx(fromRational(27400,10000000), fromRational(106700,10000000)),
		List::cons(cmplx(fromRational(-300900,10000000), fromRational(-545500,10000000)),
		List::cons(cmplx(fromRational(-756300,10000000), fromRational(543200,10000000)),
		List::cons(cmplx(fromRational(625000,10000000), fromRational(625000,10000000)),
		List::cons(cmplx(fromRational(353100,10000000), fromRational(-1029300,10000000)),
		List::cons(cmplx(fromRational(-757100,10000000), fromRational(194400,10000000)),
		List::cons(cmplx(fromRational(-441500,10000000), fromRational(665000,10000000)),
		List::cons(cmplx(fromRational(369300,10000000), fromRational(-62800,10000000)),
		List::cons(cmplx(fromRational(920500,10000000), fromRational(597200,10000000)),
		List::cons(cmplx(fromRational(347100,10000000), fromRational(-294900,10000000)),
		List::cons(cmplx(fromRational(206500,10000000), fromRational(-921400,10000000)),
		List::cons(cmplx(fromRational(552400,10000000), fromRational(-552400,10000000)),
		List::cons(cmplx(fromRational(-10100,10000000), fromRational(-169700,10000000)),
		List::cons(cmplx(fromRational(-34800,10000000), fromRational(558900,10000000)),
		List::cons(cmplx(fromRational(-239100,10000000), fromRational(-507500,10000000)),
		List::cons(cmplx(fromRational(-1021400,10000000), fromRational(-284700,10000000)),
		List::cons(cmplx(fromRational(-312000,10000000), fromRational(869900,10000000)),
		List::cons(cmplx(fromRational(766700,10000000), fromRational(-538200,10000000)),
		List::cons(cmplx(fromRational(-103800,10000000), fromRational(-519300,10000000)),
		List::cons(cmplx(fromRational(-1093800,10000000), fromRational(-156200,10000000)),
		List::cons(cmplx(fromRational(-160700,10000000), fromRational(-690600,10000000)),
		List::cons(cmplx(fromRational(-77700,10000000), fromRational(508300,10000000)),
		List::cons(cmplx(fromRational(-821800,10000000), fromRational(383000,10000000)),
		List::cons(cmplx(fromRational(-21700,10000000), fromRational(-623000,10000000)),
		List::cons(cmplx(fromRational(576500,10000000), fromRational(-112100,10000000)),
		List::cons(cmplx(fromRational(889200,10000000), fromRational(406700,10000000)),
		List::cons(cmplx(fromRational(400100,10000000), fromRational(645400,10000000)),
		List::cons(cmplx(fromRational(-773400,10000000), fromRational(773400,10000000)),
		List::cons(cmplx(fromRational(303000,10000000), fromRational(789100,10000000)),
		List::cons(cmplx(fromRational(471400,10000000), fromRational(-193200,10000000)),
		List::cons(cmplx(fromRational(-805300,10000000), fromRational(-747500,10000000)),
		List::cons(cmplx(fromRational(-359400,10000000), fromRational(753800,10000000)),
		List::cons(cmplx(fromRational(-303100,10000000), fromRational(727700,10000000)),
		List::cons(cmplx(fromRational(127500,10000000), fromRational(-13700,10000000)),
		List::cons(cmplx(fromRational(876900,10000000), fromRational(655200,10000000)),
		List::cons(cmplx(fromRational(0,10000000), fromRational(0,10000000)),
		List::cons(cmplx(fromRational(81500,10000000), fromRational(-850300,10000000)),
		List::cons(cmplx(fromRational(775300,10000000), fromRational(-753700,10000000)),
		List::cons(cmplx(fromRational(875700,10000000), fromRational(-480000,10000000)),
		List::cons(cmplx(fromRational(827100,10000000), fromRational(634200,10000000)),
		List::cons(cmplx(fromRational(328700,10000000), fromRational(629200,10000000)),
		List::cons(cmplx(fromRational(259700,10000000), fromRational(-300800,10000000)),
		List::cons(cmplx(fromRational(-244500,10000000), fromRational(337300,10000000)),
		List::cons(cmplx(fromRational(-552400,10000000), fromRational(552400,10000000)),
		List::cons(cmplx(fromRational(718800,10000000), fromRational(-143500,10000000)),
		List::cons(cmplx(fromRational(833200,10000000), fromRational(478600,10000000)),
		List::cons(cmplx(fromRational(-129400,10000000), fromRational(371600,10000000)),
		List::cons(cmplx(fromRational(83900,10000000), fromRational(-911700,10000000)),
		List::cons(cmplx(fromRational(598800,10000000), fromRational(-279400,10000000)),
		List::cons(cmplx(fromRational(214700,10000000), fromRational(655500,10000000)),
		List::cons(cmplx(fromRational(-439100,10000000), fromRational(678400,10000000)),
		List::cons(cmplx(fromRational(-781200,10000000), fromRational(781200,10000000)),
		List::cons(cmplx(fromRational(-1006600,10000000), fromRational(-149600,10000000)),
		List::cons(cmplx(fromRational(-382500,10000000), fromRational(-391000,10000000)),
		List::cons(cmplx(fromRational(-101900,10000000), fromRational(45900,10000000)),
		List::cons(cmplx(fromRational(-549600,10000000), fromRational(-573400,10000000)),
		List::cons(cmplx(fromRational(296900,10000000), fromRational(112400,10000000)),
		List::cons(cmplx(fromRational(195900,10000000), fromRational(630800,10000000)),
		List::cons(cmplx(fromRational(-306100,10000000), fromRational(-535100,10000000)),
		List::cons(cmplx(fromRational(773400,10000000), fromRational(-773400,10000000)),
		List::cons(cmplx(fromRational(87100,10000000), fromRational(-407700,10000000)),
		List::cons(cmplx(fromRational(-827800,10000000), fromRational(-402500,10000000)),
		List::cons(cmplx(fromRational(-470600,10000000), fromRational(-614400,10000000)),
		List::cons(cmplx(fromRational(-578100,10000000), fromRational(-182400,10000000)),
		List::cons(cmplx(fromRational(27400,10000000), fromRational(106700,10000000)),
		List::cons(cmplx(fromRational(-300900,10000000), fromRational(-545500,10000000)),
		List::cons(cmplx(fromRational(-756300,10000000), fromRational(543200,10000000)),
		List::cons(cmplx(fromRational(625000,10000000), fromRational(625000,10000000)),
		List::cons(cmplx(fromRational(353100,10000000), fromRational(-1029300,10000000)),
		List::cons(cmplx(fromRational(-757100,10000000), fromRational(194400,10000000)),
		List::cons(cmplx(fromRational(-441500,10000000), fromRational(665000,10000000)),
		List::cons(cmplx(fromRational(369300,10000000), fromRational(-62800,10000000)),
		List::cons(cmplx(fromRational(920500,10000000), fromRational(597200,10000000)),
		List::cons(cmplx(fromRational(347100,10000000), fromRational(-294900,10000000)),
		List::cons(cmplx(fromRational(206500,10000000), fromRational(-921400,10000000)),
		List::cons(cmplx(fromRational(552400,10000000), fromRational(-552400,10000000)),
		List::cons(cmplx(fromRational(-10100,10000000), fromRational(-169700,10000000)),
		List::cons(cmplx(fromRational(-34800,10000000), fromRational(558900,10000000)),
		List::cons(cmplx(fromRational(-239100,10000000), fromRational(-507500,10000000)),
		List::cons(cmplx(fromRational(-1021400,10000000), fromRational(-284700,10000000)),
		List::cons(cmplx(fromRational(-312000,10000000), fromRational(869900,10000000)),
		List::cons(cmplx(fromRational(766700,10000000), fromRational(-538200,10000000)),
		List::cons(cmplx(fromRational(-103800,10000000), fromRational(-519300,10000000)),
		List::cons(cmplx(fromRational(-1093800,10000000), fromRational(-156200,10000000)),
		List::cons(cmplx(fromRational(-160700,10000000), fromRational(-690600,10000000)),
		List::cons(cmplx(fromRational(-77700,10000000), fromRational(508300,10000000)),
		List::cons(cmplx(fromRational(-821800,10000000), fromRational(383000,10000000)),
		List::cons(cmplx(fromRational(-21700,10000000), fromRational(-623000,10000000)),
		List::cons(cmplx(fromRational(576500,10000000), fromRational(-112100,10000000)),
		List::cons(cmplx(fromRational(889200,10000000), fromRational(406700,10000000)),
		List::cons(cmplx(fromRational(400100,10000000), fromRational(645400,10000000)),
		List::cons(cmplx(fromRational(-773400,10000000), fromRational(773400,10000000)),
		List::cons(cmplx(fromRational(303000,10000000), fromRational(789100,10000000)),
		List::cons(cmplx(fromRational(471400,10000000), fromRational(-193200,10000000)),
		List::cons(cmplx(fromRational(-805300,10000000), fromRational(-747500,10000000)),
		List::cons(cmplx(fromRational(-359400,10000000), fromRational(753800,10000000)),
		List::cons(cmplx(fromRational(-303100,10000000), fromRational(727700,10000000)),
		List::cons(cmplx(fromRational(127500,10000000), fromRational(-13700,10000000)),
		List::cons(cmplx(fromRational(876900,10000000), fromRational(655200,10000000)),
		List::cons(cmplx(fromRational(0,10000000), fromRational(0,10000000)),
		List::cons(cmplx(fromRational(81500,10000000), fromRational(-850300,10000000)),
		List::cons(cmplx(fromRational(775300,10000000), fromRational(-753700,10000000)),
		List::cons(cmplx(fromRational(875700,10000000), fromRational(-480000,10000000)),
		List::cons(cmplx(fromRational(827100,10000000), fromRational(634200,10000000)),
		List::cons(cmplx(fromRational(328700,10000000), fromRational(629200,10000000)),
		List::cons(cmplx(fromRational(259700,10000000), fromRational(-300800,10000000)),
		List::cons(cmplx(fromRational(-244500,10000000), fromRational(337300,10000000)),
		List::cons(cmplx(fromRational(-552400,10000000), fromRational(552400,10000000)),
		List::cons(cmplx(fromRational(718800,10000000), fromRational(-143500,10000000)),
		List::cons(cmplx(fromRational(833200,10000000), fromRational(478600,10000000)),
		List::cons(cmplx(fromRational(-129400,10000000), fromRational(371600,10000000)),
		List::cons(cmplx(fromRational(83900,10000000), fromRational(-911700,10000000)),
		List::cons(cmplx(fromRational(598800,10000000), fromRational(-279400,10000000)),
		List::cons(cmplx(fromRational(214700,10000000), fromRational(655500,10000000)),
		List::cons(cmplx(fromRational(-439100,10000000), fromRational(678400,10000000)),
		List::cons(cmplx(fromRational(-781200,10000000), fromRational(781200,10000000)),
		List::cons(cmplx(fromRational(-1006600,10000000), fromRational(-149600,10000000)),
		List::cons(cmplx(fromRational(-382500,10000000), fromRational(-391000,10000000)),
		List::cons(cmplx(fromRational(-101900,10000000), fromRational(45900,10000000)),
		List::cons(cmplx(fromRational(-549600,10000000), fromRational(-573400,10000000)),
		List::cons(cmplx(fromRational(296900,10000000), fromRational(112400,10000000)),
		List::cons(cmplx(fromRational(195900,10000000), fromRational(630800,10000000)),
		List::cons(cmplx(fromRational(-306100,10000000), fromRational(-535100,10000000)),
		List::cons(cmplx(fromRational(773400,10000000), fromRational(-773400,10000000)),
		List::cons(cmplx(fromRational(87100,10000000), fromRational(-407700,10000000)),
		List::cons(cmplx(fromRational(-827800,10000000), fromRational(-402500,10000000)),
		List::cons(cmplx(fromRational(-470600,10000000), fromRational(-614400,10000000)),
		List::cons(cmplx(fromRational(-578100,10000000), fromRational(-182400,10000000)),
		List::cons(cmplx(fromRational(27400,10000000), fromRational(106700,10000000)),
		List::cons(cmplx(fromRational(-300900,10000000), fromRational(-545500,10000000)),
		List::cons(cmplx(fromRational(-756300,10000000), fromRational(543200,10000000)),
		List::nil)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
	return tempV;
endfunction

// function to generate long training sequence
function Vector#(256, FPComplex#(2,14)) getLongPreambles();
	Vector#(256, FPComplex#(2,14)) tempV = Vector::toVector(
		List::cons(cmplx(fromRational(441900,10000000), fromRational(441900,10000000)),
		List::cons(cmplx(fromRational(865600,10000000), fromRational(-503600,10000000)),
		List::cons(cmplx(fromRational(-626200,10000000), fromRational(31200,10000000)),
		List::cons(cmplx(fromRational(-689100,10000000), fromRational(-100900,10000000)),
		List::cons(cmplx(fromRational(573600,10000000), fromRational(-273000,10000000)),
		List::cons(cmplx(fromRational(466500,10000000), fromRational(843300,10000000)),
		List::cons(cmplx(fromRational(-335900,10000000), fromRational(-59200,10000000)),
		List::cons(cmplx(fromRational(271400,10000000), fromRational(-1032800,10000000)),
		List::cons(cmplx(fromRational(890700,10000000), fromRational(-467900,10000000)),
		List::cons(cmplx(fromRational(641400,10000000), fromRational(92200,10000000)),
		List::cons(cmplx(fromRational(553600,10000000), fromRational(840900,10000000)),
		List::cons(cmplx(fromRational(-388100,10000000), fromRational(245800,10000000)),
		List::cons(cmplx(fromRational(-919600,10000000), fromRational(219300,10000000)),
		List::cons(cmplx(fromRational(167900,10000000), fromRational(1029600,10000000)),
		List::cons(cmplx(fromRational(339600,10000000), fromRational(-565000,10000000)),
		List::cons(cmplx(fromRational(-453400,10000000), fromRational(-756300,10000000)),
		List::cons(cmplx(fromRational(-851500,10000000), fromRational(436400,10000000)),
		List::cons(cmplx(fromRational(-718100,10000000), fromRational(-66900,10000000)),
		List::cons(cmplx(fromRational(-281400,10000000), fromRational(577000,10000000)),
		List::cons(cmplx(fromRational(-226800,10000000), fromRational(953700,10000000)),
		List::cons(cmplx(fromRational(-144900,10000000), fromRational(-75600,10000000)),
		List::cons(cmplx(fromRational(357800,10000000), fromRational(-65900,10000000)),
		List::cons(cmplx(fromRational(880600,10000000), fromRational(-134900,10000000)),
		List::cons(cmplx(fromRational(575500,10000000), fromRational(111600,10000000)),
		List::cons(cmplx(fromRational(-36500,10000000), fromRational(1057300,10000000)),
		List::cons(cmplx(fromRational(760700,10000000), fromRational(539600,10000000)),
		List::cons(cmplx(fromRational(589000,10000000), fromRational(-453000,10000000)),
		List::cons(cmplx(fromRational(-1002600,10000000), fromRational(-127200,10000000)),
		List::cons(cmplx(fromRational(-390000,10000000), fromRational(636700,10000000)),
		List::cons(cmplx(fromRational(450300,10000000), fromRational(778700,10000000)),
		List::cons(cmplx(fromRational(123400,10000000), fromRational(729700,10000000)),
		List::cons(cmplx(fromRational(713300,10000000), fromRational(503300,10000000)),
		List::cons(cmplx(fromRational(773400,10000000), fromRational(-110500,10000000)),
		List::cons(cmplx(fromRational(398400,10000000), fromRational(-230700,10000000)),
		List::cons(cmplx(fromRational(622200,10000000), fromRational(-413600,10000000)),
		List::cons(cmplx(fromRational(277500,10000000), fromRational(-560600,10000000)),
		List::cons(cmplx(fromRational(456700,10000000), fromRational(334600,10000000)),
		List::cons(cmplx(fromRational(833700,10000000), fromRational(-4900,10000000)),
		List::cons(cmplx(fromRational(-155100,10000000), fromRational(-872800,10000000)),
		List::cons(cmplx(fromRational(-468800,10000000), fromRational(557000,10000000)),
		List::cons(cmplx(fromRational(239300,10000000), fromRational(781400,10000000)),
		List::cons(cmplx(fromRational(601800,10000000), fromRational(-765600,10000000)),
		List::cons(cmplx(fromRational(707800,10000000), fromRational(-158200,10000000)),
		List::cons(cmplx(fromRational(-240000,10000000), fromRational(253200,10000000)),
		List::cons(cmplx(fromRational(-716200,10000000), fromRational(-660000,10000000)),
		List::cons(cmplx(fromRational(410400,10000000), fromRational(-71200,10000000)),
		List::cons(cmplx(fromRational(363400,10000000), fromRational(847700,10000000)),
		List::cons(cmplx(fromRational(-100300,10000000), fromRational(1094700,10000000)),
		List::cons(cmplx(fromRational(-318100,10000000), fromRational(786800,10000000)),
		List::cons(cmplx(fromRational(-1031000,10000000), fromRational(174100,10000000)),
		List::cons(cmplx(fromRational(107500,10000000), fromRational(272800,10000000)),
		List::cons(cmplx(fromRational(533600,10000000), fromRational(-432600,10000000)),
		List::cons(cmplx(fromRational(-873800,10000000), fromRational(-670400,10000000)),
		List::cons(cmplx(fromRational(-55900,10000000), fromRational(782700,10000000)),
		List::cons(cmplx(fromRational(713000,10000000), fromRational(495700,10000000)),
		List::cons(cmplx(fromRational(478900,10000000), fromRational(-294300,10000000)),
		List::cons(cmplx(fromRational(758300,10000000), fromRational(-335500,10000000)),
		List::cons(cmplx(fromRational(22300,10000000), fromRational(-955800,10000000)),
		List::cons(cmplx(fromRational(-128900,10000000), fromRational(-609300,10000000)),
		List::cons(cmplx(fromRational(60500,10000000), fromRational(-49600,10000000)),
		List::cons(cmplx(fromRational(-389100,10000000), fromRational(482200,10000000)),
		List::cons(cmplx(fromRational(-260300,10000000), fromRational(796600,10000000)),
		List::cons(cmplx(fromRational(-907700,10000000), fromRational(-165000,10000000)),
		List::cons(cmplx(fromRational(-667400,10000000), fromRational(374500,10000000)),
		List::cons(cmplx(fromRational(441900,10000000), fromRational(441900,10000000)),
		List::cons(cmplx(fromRational(-366300,10000000), fromRational(-952100,10000000)),
		List::cons(cmplx(fromRational(-444600,10000000), fromRational(243800,10000000)),
		List::cons(cmplx(fromRational(64800,10000000), fromRational(1041400,10000000)),
		List::cons(cmplx(fromRational(-51300,10000000), fromRational(184200,10000000)),
		List::cons(cmplx(fromRational(835400,10000000), fromRational(1300,10000000)),
		List::cons(cmplx(fromRational(826800,10000000), fromRational(-357800,10000000)),
		List::cons(cmplx(fromRational(20600,10000000), fromRational(-270300,10000000)),
		List::cons(cmplx(fromRational(-109500,10000000), fromRational(-313300,10000000)),
		List::cons(cmplx(fromRational(-655700,10000000), fromRational(-332100,10000000)),
		List::cons(cmplx(fromRational(-602900,10000000), fromRational(-50400,10000000)),
		List::cons(cmplx(fromRational(49900,10000000), fromRational(-963600,10000000)),
		List::cons(cmplx(fromRational(-524900,10000000), fromRational(-622000,10000000)),
		List::cons(cmplx(fromRational(-609100,10000000), fromRational(200600,10000000)),
		List::cons(cmplx(fromRational(744800,10000000), fromRational(-196100,10000000)),
		List::cons(cmplx(fromRational(306700,10000000), fromRational(21900,10000000)),
		List::cons(cmplx(fromRational(-695300,10000000), fromRational(-657400,10000000)),
		List::cons(cmplx(fromRational(490900,10000000), fromRational(-909800,10000000)),
		List::cons(cmplx(fromRational(171600,10000000), fromRational(141800,10000000)),
		List::cons(cmplx(fromRational(-935400,10000000), fromRational(-412100,10000000)),
		List::cons(cmplx(fromRational(114100,10000000), fromRational(-805400,10000000)),
		List::cons(cmplx(fromRational(457500,10000000), fromRational(-92600,10000000)),
		List::cons(cmplx(fromRational(377000,10000000), fromRational(710100,10000000)),
		List::cons(cmplx(fromRational(-9600,10000000), fromRational(801200,10000000)),
		List::cons(cmplx(fromRational(-1057300,10000000), fromRational(36500,10000000)),
		List::cons(cmplx(fromRational(-332200,10000000), fromRational(576300,10000000)),
		List::cons(cmplx(fromRational(77600,10000000), fromRational(179900,10000000)),
		List::cons(cmplx(fromRational(-136300,10000000), fromRational(-929900,10000000)),
		List::cons(cmplx(fromRational(-118300,10000000), fromRational(429300,10000000)),
		List::cons(cmplx(fromRational(-878900,10000000), fromRational(250400,10000000)),
		List::cons(cmplx(fromRational(56900,10000000), fromRational(-749100,10000000)),
		List::cons(cmplx(fromRational(526900,10000000), fromRational(423300,10000000)),
		List::cons(cmplx(fromRational(-773400,10000000), fromRational(110500,10000000)),
		List::cons(cmplx(fromRational(-283100,10000000), fromRational(-971700,10000000)),
		List::cons(cmplx(fromRational(474300,10000000), fromRational(-652300,10000000)),
		List::cons(cmplx(fromRational(960900,10000000), fromRational(-118300,10000000)),
		List::cons(cmplx(fromRational(713000,10000000), fromRational(562300,10000000)),
		List::cons(cmplx(fromRational(-368800,10000000), fromRational(894700,10000000)),
		List::cons(cmplx(fromRational(522300,10000000), fromRational(447400,10000000)),
		List::cons(cmplx(fromRational(123100,10000000), fromRational(-79900,10000000)),
		List::cons(cmplx(fromRational(-1020600,10000000), fromRational(-200,10000000)),
		List::cons(cmplx(fromRational(414700,10000000), fromRational(562700,10000000)),
		List::cons(cmplx(fromRational(470600,10000000), fromRational(835100,10000000)),
		List::cons(cmplx(fromRational(57000,10000000), fromRational(272400,10000000)),
		List::cons(cmplx(fromRational(834800,10000000), fromRational(-629300,10000000)),
		List::cons(cmplx(fromRational(436400,10000000), fromRational(-323900,10000000)),
		List::cons(cmplx(fromRational(-59800,10000000), fromRational(79200,10000000)),
		List::cons(cmplx(fromRational(-520700,10000000), fromRational(-135300,10000000)),
		List::cons(cmplx(fromRational(-786800,10000000), fromRational(318100,10000000)),
		List::cons(cmplx(fromRational(-392500,10000000), fromRational(-385700,10000000)),
		List::cons(cmplx(fromRational(-648400,10000000), fromRational(-825800,10000000)),
		List::cons(cmplx(fromRational(-677800,10000000), fromRational(497400,10000000)),
		List::cons(cmplx(fromRational(96500,10000000), fromRational(-140600,10000000)),
		List::cons(cmplx(fromRational(475800,10000000), fromRational(-623700,10000000)),
		List::cons(cmplx(fromRational(-435900,10000000), fromRational(396400,10000000)),
		List::cons(cmplx(fromRational(-911800,10000000), fromRational(-462500,10000000)),
		List::cons(cmplx(fromRational(335500,10000000), fromRational(-758300,10000000)),
		List::cons(cmplx(fromRational(100900,10000000), fromRational(379200,10000000)),
		List::cons(cmplx(fromRational(-1041800,10000000), fromRational(40100,10000000)),
		List::cons(cmplx(fromRational(-726000,10000000), fromRational(-819300,10000000)),
		List::cons(cmplx(fromRational(-428400,10000000), fromRational(-740200,10000000)),
		List::cons(cmplx(fromRational(299100,10000000), fromRational(-645700,10000000)),
		List::cons(cmplx(fromRational(482200,10000000), fromRational(-606400,10000000)),
		List::cons(cmplx(fromRational(-402200,10000000), fromRational(393800,10000000)),
		List::cons(cmplx(fromRational(441900,10000000), fromRational(441900,10000000)),
		List::cons(cmplx(fromRational(865600,10000000), fromRational(-503600,10000000)),
		List::cons(cmplx(fromRational(-626200,10000000), fromRational(31200,10000000)),
		List::cons(cmplx(fromRational(-689100,10000000), fromRational(-100900,10000000)),
		List::cons(cmplx(fromRational(573600,10000000), fromRational(-273000,10000000)),
		List::cons(cmplx(fromRational(466500,10000000), fromRational(843300,10000000)),
		List::cons(cmplx(fromRational(-335900,10000000), fromRational(-59200,10000000)),
		List::cons(cmplx(fromRational(271400,10000000), fromRational(-1032800,10000000)),
		List::cons(cmplx(fromRational(890700,10000000), fromRational(-467900,10000000)),
		List::cons(cmplx(fromRational(641400,10000000), fromRational(92200,10000000)),
		List::cons(cmplx(fromRational(553600,10000000), fromRational(840900,10000000)),
		List::cons(cmplx(fromRational(-388100,10000000), fromRational(245800,10000000)),
		List::cons(cmplx(fromRational(-919600,10000000), fromRational(219300,10000000)),
		List::cons(cmplx(fromRational(167900,10000000), fromRational(1029600,10000000)),
		List::cons(cmplx(fromRational(339600,10000000), fromRational(-565000,10000000)),
		List::cons(cmplx(fromRational(-453400,10000000), fromRational(-756300,10000000)),
		List::cons(cmplx(fromRational(-851500,10000000), fromRational(436400,10000000)),
		List::cons(cmplx(fromRational(-718100,10000000), fromRational(-66900,10000000)),
		List::cons(cmplx(fromRational(-281400,10000000), fromRational(577000,10000000)),
		List::cons(cmplx(fromRational(-226800,10000000), fromRational(953700,10000000)),
		List::cons(cmplx(fromRational(-144900,10000000), fromRational(-75600,10000000)),
		List::cons(cmplx(fromRational(357800,10000000), fromRational(-65900,10000000)),
		List::cons(cmplx(fromRational(880600,10000000), fromRational(-134900,10000000)),
		List::cons(cmplx(fromRational(575500,10000000), fromRational(111600,10000000)),
		List::cons(cmplx(fromRational(-36500,10000000), fromRational(1057300,10000000)),
		List::cons(cmplx(fromRational(760700,10000000), fromRational(539600,10000000)),
		List::cons(cmplx(fromRational(589000,10000000), fromRational(-453000,10000000)),
		List::cons(cmplx(fromRational(-1002600,10000000), fromRational(-127200,10000000)),
		List::cons(cmplx(fromRational(-390000,10000000), fromRational(636700,10000000)),
		List::cons(cmplx(fromRational(450300,10000000), fromRational(778700,10000000)),
		List::cons(cmplx(fromRational(123400,10000000), fromRational(729700,10000000)),
		List::cons(cmplx(fromRational(713300,10000000), fromRational(503300,10000000)),
		List::cons(cmplx(fromRational(773400,10000000), fromRational(-110500,10000000)),
		List::cons(cmplx(fromRational(398400,10000000), fromRational(-230700,10000000)),
		List::cons(cmplx(fromRational(622200,10000000), fromRational(-413600,10000000)),
		List::cons(cmplx(fromRational(277500,10000000), fromRational(-560600,10000000)),
		List::cons(cmplx(fromRational(456700,10000000), fromRational(334600,10000000)),
		List::cons(cmplx(fromRational(833700,10000000), fromRational(-4900,10000000)),
		List::cons(cmplx(fromRational(-155100,10000000), fromRational(-872800,10000000)),
		List::cons(cmplx(fromRational(-468800,10000000), fromRational(557000,10000000)),
		List::cons(cmplx(fromRational(239300,10000000), fromRational(781400,10000000)),
		List::cons(cmplx(fromRational(601800,10000000), fromRational(-765600,10000000)),
		List::cons(cmplx(fromRational(707800,10000000), fromRational(-158200,10000000)),
		List::cons(cmplx(fromRational(-240000,10000000), fromRational(253200,10000000)),
		List::cons(cmplx(fromRational(-716200,10000000), fromRational(-660000,10000000)),
		List::cons(cmplx(fromRational(410400,10000000), fromRational(-71200,10000000)),
		List::cons(cmplx(fromRational(363400,10000000), fromRational(847700,10000000)),
		List::cons(cmplx(fromRational(-100300,10000000), fromRational(1094700,10000000)),
		List::cons(cmplx(fromRational(-318100,10000000), fromRational(786800,10000000)),
		List::cons(cmplx(fromRational(-1031000,10000000), fromRational(174100,10000000)),
		List::cons(cmplx(fromRational(107500,10000000), fromRational(272800,10000000)),
		List::cons(cmplx(fromRational(533600,10000000), fromRational(-432600,10000000)),
		List::cons(cmplx(fromRational(-873800,10000000), fromRational(-670400,10000000)),
		List::cons(cmplx(fromRational(-55900,10000000), fromRational(782700,10000000)),
		List::cons(cmplx(fromRational(713000,10000000), fromRational(495700,10000000)),
		List::cons(cmplx(fromRational(478900,10000000), fromRational(-294300,10000000)),
		List::cons(cmplx(fromRational(758300,10000000), fromRational(-335500,10000000)),
		List::cons(cmplx(fromRational(22300,10000000), fromRational(-955800,10000000)),
		List::cons(cmplx(fromRational(-128900,10000000), fromRational(-609300,10000000)),
		List::cons(cmplx(fromRational(60500,10000000), fromRational(-49600,10000000)),
		List::cons(cmplx(fromRational(-389100,10000000), fromRational(482200,10000000)),
		List::cons(cmplx(fromRational(-260300,10000000), fromRational(796600,10000000)),
		List::cons(cmplx(fromRational(-907700,10000000), fromRational(-165000,10000000)),
		List::cons(cmplx(fromRational(-667400,10000000), fromRational(374500,10000000)),
		List::cons(cmplx(fromRational(441900,10000000), fromRational(441900,10000000)),
		List::cons(cmplx(fromRational(-366300,10000000), fromRational(-952100,10000000)),
		List::cons(cmplx(fromRational(-444600,10000000), fromRational(243800,10000000)),
		List::cons(cmplx(fromRational(64800,10000000), fromRational(1041400,10000000)),
		List::cons(cmplx(fromRational(-51300,10000000), fromRational(184200,10000000)),
		List::cons(cmplx(fromRational(835400,10000000), fromRational(1300,10000000)),
		List::cons(cmplx(fromRational(826800,10000000), fromRational(-357800,10000000)),
		List::cons(cmplx(fromRational(20600,10000000), fromRational(-270300,10000000)),
		List::cons(cmplx(fromRational(-109500,10000000), fromRational(-313300,10000000)),
		List::cons(cmplx(fromRational(-655700,10000000), fromRational(-332100,10000000)),
		List::cons(cmplx(fromRational(-602900,10000000), fromRational(-50400,10000000)),
		List::cons(cmplx(fromRational(49900,10000000), fromRational(-963600,10000000)),
		List::cons(cmplx(fromRational(-524900,10000000), fromRational(-622000,10000000)),
		List::cons(cmplx(fromRational(-609100,10000000), fromRational(200600,10000000)),
		List::cons(cmplx(fromRational(744800,10000000), fromRational(-196100,10000000)),
		List::cons(cmplx(fromRational(306700,10000000), fromRational(21900,10000000)),
		List::cons(cmplx(fromRational(-695300,10000000), fromRational(-657400,10000000)),
		List::cons(cmplx(fromRational(490900,10000000), fromRational(-909800,10000000)),
		List::cons(cmplx(fromRational(171600,10000000), fromRational(141800,10000000)),
		List::cons(cmplx(fromRational(-935400,10000000), fromRational(-412100,10000000)),
		List::cons(cmplx(fromRational(114100,10000000), fromRational(-805400,10000000)),
		List::cons(cmplx(fromRational(457500,10000000), fromRational(-92600,10000000)),
		List::cons(cmplx(fromRational(377000,10000000), fromRational(710100,10000000)),
		List::cons(cmplx(fromRational(-9600,10000000), fromRational(801200,10000000)),
		List::cons(cmplx(fromRational(-1057300,10000000), fromRational(36500,10000000)),
		List::cons(cmplx(fromRational(-332200,10000000), fromRational(576300,10000000)),
		List::cons(cmplx(fromRational(77600,10000000), fromRational(179900,10000000)),
		List::cons(cmplx(fromRational(-136300,10000000), fromRational(-929900,10000000)),
		List::cons(cmplx(fromRational(-118300,10000000), fromRational(429300,10000000)),
		List::cons(cmplx(fromRational(-878900,10000000), fromRational(250400,10000000)),
		List::cons(cmplx(fromRational(56900,10000000), fromRational(-749100,10000000)),
		List::cons(cmplx(fromRational(526900,10000000), fromRational(423300,10000000)),
		List::cons(cmplx(fromRational(-773400,10000000), fromRational(110500,10000000)),
		List::cons(cmplx(fromRational(-283100,10000000), fromRational(-971700,10000000)),
		List::cons(cmplx(fromRational(474300,10000000), fromRational(-652300,10000000)),
		List::cons(cmplx(fromRational(960900,10000000), fromRational(-118300,10000000)),
		List::cons(cmplx(fromRational(713000,10000000), fromRational(562300,10000000)),
		List::cons(cmplx(fromRational(-368800,10000000), fromRational(894700,10000000)),
		List::cons(cmplx(fromRational(522300,10000000), fromRational(447400,10000000)),
		List::cons(cmplx(fromRational(123100,10000000), fromRational(-79900,10000000)),
		List::cons(cmplx(fromRational(-1020600,10000000), fromRational(-200,10000000)),
		List::cons(cmplx(fromRational(414700,10000000), fromRational(562700,10000000)),
		List::cons(cmplx(fromRational(470600,10000000), fromRational(835100,10000000)),
		List::cons(cmplx(fromRational(57000,10000000), fromRational(272400,10000000)),
		List::cons(cmplx(fromRational(834800,10000000), fromRational(-629300,10000000)),
		List::cons(cmplx(fromRational(436400,10000000), fromRational(-323900,10000000)),
		List::cons(cmplx(fromRational(-59800,10000000), fromRational(79200,10000000)),
		List::cons(cmplx(fromRational(-520700,10000000), fromRational(-135300,10000000)),
		List::cons(cmplx(fromRational(-786800,10000000), fromRational(318100,10000000)),
		List::cons(cmplx(fromRational(-392500,10000000), fromRational(-385700,10000000)),
		List::cons(cmplx(fromRational(-648400,10000000), fromRational(-825800,10000000)),
		List::cons(cmplx(fromRational(-677800,10000000), fromRational(497400,10000000)),
		List::cons(cmplx(fromRational(96500,10000000), fromRational(-140600,10000000)),
		List::cons(cmplx(fromRational(475800,10000000), fromRational(-623700,10000000)),
		List::cons(cmplx(fromRational(-435900,10000000), fromRational(396400,10000000)),
		List::cons(cmplx(fromRational(-911800,10000000), fromRational(-462500,10000000)),
		List::cons(cmplx(fromRational(335500,10000000), fromRational(-758300,10000000)),
		List::cons(cmplx(fromRational(100900,10000000), fromRational(379200,10000000)),
		List::cons(cmplx(fromRational(-1041800,10000000), fromRational(40100,10000000)),
		List::cons(cmplx(fromRational(-726000,10000000), fromRational(-819300,10000000)),
		List::cons(cmplx(fromRational(-428400,10000000), fromRational(-740200,10000000)),
		List::cons(cmplx(fromRational(299100,10000000), fromRational(-645700,10000000)),
		List::cons(cmplx(fromRational(482200,10000000), fromRational(-606400,10000000)),
		List::cons(cmplx(fromRational(-402200,10000000), fromRational(393800,10000000)),
		List::nil)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
	return tempV;
endfunction

// function to generate long training sequence (signs only)
function Vector#(256, Complex#(Bit#(1))) getLongPreSigns();
	Vector#(256, Complex#(Bit#(1))) tempV = Vector::toVector(
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 0),
		List::cons(cmplx(1, 0),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(1, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(0, 1),
		List::cons(cmplx(1, 0),
		List::nil)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
	return tempV;
endfunction

// module to generate sample packet
(* synthesize *)
module mkPacket(RegFile#(Bit#(10), FPComplex#(2,14)));
	RegFile#(Bit#(10), FPComplex#(2,14)) regFile <- mkRegFileLoad("WiMAXPacket.txt",0,1023);
	return regFile;
endmodule

// module to generate sample packet
(* synthesize *)
module mkTweakedPacket(RegFile#(Bit#(10), FPComplex#(2,14)));
	RegFile#(Bit#(10), FPComplex#(2,14)) regFile <- mkRegFileLoad("WiMAXTweakedPacket.txt",0,1023);
	return regFile;
endmodule

